** Profile: "SCHEMATIC1-Switch sim profile"  [ C:\USERS\MATTHEW EINHORN\DESKTOP\CPL ADC BOARD\Boutput board\Simulation\switch sim-pspicefiles\schematic1\switch sim profile.sim ] 

** Creating circuit file "Switch sim profile.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "C:\USERS\MATTHEW EINHORN\DESKTOP\CPL ADC BOARD\Boutput board\Simulation\switch sim-pspicefiles\schematic1\Switch sim profile\"
+ "Switch sim profile_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Matthew Einhorn\Documents\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 3.0001 2 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
